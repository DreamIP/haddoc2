library ieee;
	use	ieee.std_logic_1164.all;

end package cnn_kernels is
    
end package;
